module bitonicMerge #(

)(

)

endmodule